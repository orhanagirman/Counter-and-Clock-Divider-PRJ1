----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:57:53 08/03/2020 
-- Design Name: 
-- Module Name:    three_bit_bicounter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity three_bit_bicounter is
    Port ( clk : in STD_LOGIC;
	        rst : in  STD_LOGIC;
           x : in  STD_LOGIC;
           output : out  STD_LOGIC_VECTOR (2 downto 0));
end three_bit_bicounter;

architecture Behavioral of three_bit_bicounter is
Signal count: STD_LOGIC_VECTOR (2 downto 0);

begin
   process(rst,clk)
   begin
      if (rst = '1') then
          count <= "000";
      elsif (clk'EVENT) and (clk = '1') then
             if (x = '1') then
                 count <= count + 1;
				 elsif (x = '0') then
                 count <= count - 1;				 
             end if;
	   end if;	
	end process;	
	output <= count;




end Behavioral;

